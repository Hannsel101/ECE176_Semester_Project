module RegisterFile(
	input [2:0] R1, R2, R3,//Register pointers
	input [12:0] ALU_Result,//Result from the ALU arithmetic operation
	input WriteFlag);//Flag to enable a write into a register
	
	
	
endmodule
